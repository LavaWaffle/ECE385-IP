
module ece385_not(
    input logic op,
    output logic res
    );
    assign res = ~op;
endmodule